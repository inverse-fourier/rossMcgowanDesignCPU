`ifndef DEFS_SV
`define DEFS_SV

// Data width for registers and bus 
`define DATA_WIDTH 16

// Address width for RAM (256 bytes = 8-bit address)
`define ADDR_WIDTH 16

`endif
